//  A testbench for SumadorRestador_tb
`timescale 1us/1ns

module SumadorRestador_tb;
    reg B3;
    reg A0;
    reg A1;
    reg A2;
    reg A3;
    reg B2;
    reg B1;
    reg B0;
    wire S3;
    wire S2;
    wire S1;
    wire S0;

  SumadorRestador SumadorRestador0 (
    .B3(B3),
    .A0(A0),
    .A1(A1),
    .A2(A2),
    .A3(A3),
    .B2(B2),
    .B1(B1),
    .B0(B0),
    .S3(S3),
    .S2(S2),
    .S1(S1),
    .S0(S0)
  );

    reg [11:0] patterns[0:255];
    integer i;

    initial begin
      patterns[0] = 12'b0_0_0_0_0_0_0_0_0_0_0_0;
      patterns[1] = 12'b0_0_0_0_0_0_0_1_0_0_0_1;
      patterns[2] = 12'b0_0_0_0_0_0_1_0_0_0_1_0;
      patterns[3] = 12'b0_0_0_0_0_0_1_1_0_0_1_1;
      patterns[4] = 12'b0_0_0_0_0_1_0_0_0_1_0_0;
      patterns[5] = 12'b0_0_0_0_0_1_0_1_0_1_0_1;
      patterns[6] = 12'b0_0_0_0_0_1_1_0_0_1_1_0;
      patterns[7] = 12'b0_0_0_0_0_1_1_1_0_1_1_1;
      patterns[8] = 12'b0_0_0_0_1_0_0_0_1_0_0_0;
      patterns[9] = 12'b0_0_0_0_1_0_0_1_0_1_1_1;
      patterns[10] = 12'b0_0_0_0_1_0_1_0_0_1_1_0;
      patterns[11] = 12'b0_0_0_0_1_0_1_1_0_1_0_1;
      patterns[12] = 12'b0_0_0_0_1_1_0_0_0_1_0_0;
      patterns[13] = 12'b0_0_0_0_1_1_0_1_0_0_1_1;
      patterns[14] = 12'b0_0_0_0_1_1_1_0_0_0_1_0;
      patterns[15] = 12'b0_0_0_0_1_1_1_1_0_0_0_1;
      patterns[16] = 12'b0_0_0_1_0_0_0_0_0_1_0_0;
      patterns[17] = 12'b0_0_0_1_0_0_0_1_0_0_1_1;
      patterns[18] = 12'b0_0_0_1_0_0_1_0_0_0_1_0;
      patterns[19] = 12'b0_0_0_1_0_0_1_1_0_0_0_1;
      patterns[20] = 12'b0_0_0_1_0_1_0_0_0_0_0_0;
      patterns[21] = 12'b0_0_0_1_0_1_0_1_0_0_0_1;
      patterns[22] = 12'b0_0_0_1_0_1_1_0_0_0_1_0;
      patterns[23] = 12'b0_0_0_1_0_1_1_1_0_0_1_1;
      patterns[24] = 12'b0_0_0_1_1_0_0_0_1_1_0_0;
      patterns[25] = 12'b0_0_0_1_1_0_0_1_1_0_1_1;
      patterns[26] = 12'b0_0_0_1_1_0_1_0_1_0_1_0;
      patterns[27] = 12'b0_0_0_1_1_0_1_1_1_0_0_1;
      patterns[28] = 12'b0_0_0_1_1_1_0_0_1_0_0_0;
      patterns[29] = 12'b0_0_0_1_1_1_0_1_0_1_1_1;
      patterns[30] = 12'b0_0_0_1_1_1_1_0_0_1_1_0;
      patterns[31] = 12'b0_0_0_1_1_1_1_1_0_1_0_1;
      patterns[32] = 12'b0_0_1_0_0_0_0_0_0_0_1_0;
      patterns[33] = 12'b0_0_1_0_0_0_0_1_0_0_0_1;
      patterns[34] = 12'b0_0_1_0_0_0_1_0_0_0_0_0;
      patterns[35] = 12'b0_0_1_0_0_0_1_1_0_0_0_1;
      patterns[36] = 12'b0_0_1_0_0_1_0_0_0_0_1_0;
      patterns[37] = 12'b0_0_1_0_0_1_0_1_0_0_1_1;
      patterns[38] = 12'b0_0_1_0_0_1_1_0_0_1_0_0;
      patterns[39] = 12'b0_0_1_0_0_1_1_1_0_1_0_1;
      patterns[40] = 12'b0_0_1_0_1_0_0_0_1_0_1_0;
      patterns[41] = 12'b0_0_1_0_1_0_0_1_1_0_0_1;
      patterns[42] = 12'b0_0_1_0_1_0_1_0_1_0_0_0;
      patterns[43] = 12'b0_0_1_0_1_0_1_1_0_1_1_1;
      patterns[44] = 12'b0_0_1_0_1_1_0_0_0_1_1_0;
      patterns[45] = 12'b0_0_1_0_1_1_0_1_0_1_0_1;
      patterns[46] = 12'b0_0_1_0_1_1_1_0_0_1_0_0;
      patterns[47] = 12'b0_0_1_0_1_1_1_1_0_0_1_1;
      patterns[48] = 12'b0_0_1_1_0_0_0_0_0_1_1_0;
      patterns[49] = 12'b0_0_1_1_0_0_0_1_0_1_0_1;
      patterns[50] = 12'b0_0_1_1_0_0_1_0_0_1_0_0;
      patterns[51] = 12'b0_0_1_1_0_0_1_1_0_0_1_1;
      patterns[52] = 12'b0_0_1_1_0_1_0_0_0_0_1_0;
      patterns[53] = 12'b0_0_1_1_0_1_0_1_0_0_0_1;
      patterns[54] = 12'b0_0_1_1_0_1_1_0_0_0_0_0;
      patterns[55] = 12'b0_0_1_1_0_1_1_1_0_0_0_1;
      patterns[56] = 12'b0_0_1_1_1_0_0_0_1_1_1_0;
      patterns[57] = 12'b0_0_1_1_1_0_0_1_1_1_0_1;
      patterns[58] = 12'b0_0_1_1_1_0_1_0_1_1_0_0;
      patterns[59] = 12'b0_0_1_1_1_0_1_1_1_0_1_1;
      patterns[60] = 12'b0_0_1_1_1_1_0_0_1_0_1_0;
      patterns[61] = 12'b0_0_1_1_1_1_0_1_1_0_0_1;
      patterns[62] = 12'b0_0_1_1_1_1_1_0_1_0_0_0;
      patterns[63] = 12'b0_0_1_1_1_1_1_1_0_1_1_1;
      patterns[64] = 12'b0_1_0_0_0_0_0_0_0_0_0_1;
      patterns[65] = 12'b0_1_0_0_0_0_0_1_0_0_0_0;
      patterns[66] = 12'b0_1_0_0_0_0_1_0_0_0_0_1;
      patterns[67] = 12'b0_1_0_0_0_0_1_1_0_0_1_0;
      patterns[68] = 12'b0_1_0_0_0_1_0_0_0_0_1_1;
      patterns[69] = 12'b0_1_0_0_0_1_0_1_0_1_0_0;
      patterns[70] = 12'b0_1_0_0_0_1_1_0_0_1_0_1;
      patterns[71] = 12'b0_1_0_0_0_1_1_1_0_1_1_0;
      patterns[72] = 12'b0_1_0_0_1_0_0_0_1_0_0_1;
      patterns[73] = 12'b0_1_0_0_1_0_0_1_1_0_0_0;
      patterns[74] = 12'b0_1_0_0_1_0_1_0_0_1_1_1;
      patterns[75] = 12'b0_1_0_0_1_0_1_1_0_1_1_0;
      patterns[76] = 12'b0_1_0_0_1_1_0_0_0_1_0_1;
      patterns[77] = 12'b0_1_0_0_1_1_0_1_0_1_0_0;
      patterns[78] = 12'b0_1_0_0_1_1_1_0_0_0_1_1;
      patterns[79] = 12'b0_1_0_0_1_1_1_1_0_0_1_0;
      patterns[80] = 12'b0_1_0_1_0_0_0_0_0_1_0_1;
      patterns[81] = 12'b0_1_0_1_0_0_0_1_0_1_0_0;
      patterns[82] = 12'b0_1_0_1_0_0_1_0_0_0_1_1;
      patterns[83] = 12'b0_1_0_1_0_0_1_1_0_0_1_0;
      patterns[84] = 12'b0_1_0_1_0_1_0_0_0_0_0_1;
      patterns[85] = 12'b0_1_0_1_0_1_0_1_0_0_0_0;
      patterns[86] = 12'b0_1_0_1_0_1_1_0_0_0_0_1;
      patterns[87] = 12'b0_1_0_1_0_1_1_1_0_0_1_0;
      patterns[88] = 12'b0_1_0_1_1_0_0_0_1_1_0_1;
      patterns[89] = 12'b0_1_0_1_1_0_0_1_1_1_0_0;
      patterns[90] = 12'b0_1_0_1_1_0_1_0_1_0_1_1;
      patterns[91] = 12'b0_1_0_1_1_0_1_1_1_0_1_0;
      patterns[92] = 12'b0_1_0_1_1_1_0_0_1_0_0_1;
      patterns[93] = 12'b0_1_0_1_1_1_0_1_1_0_0_0;
      patterns[94] = 12'b0_1_0_1_1_1_1_0_0_1_1_1;
      patterns[95] = 12'b0_1_0_1_1_1_1_1_0_1_1_0;
      patterns[96] = 12'b0_1_1_0_0_0_0_0_0_0_1_1;
      patterns[97] = 12'b0_1_1_0_0_0_0_1_0_0_1_0;
      patterns[98] = 12'b0_1_1_0_0_0_1_0_0_0_0_1;
      patterns[99] = 12'b0_1_1_0_0_0_1_1_0_0_0_0;
      patterns[100] = 12'b0_1_1_0_0_1_0_0_0_0_0_1;
      patterns[101] = 12'b0_1_1_0_0_1_0_1_0_0_1_0;
      patterns[102] = 12'b0_1_1_0_0_1_1_0_0_0_1_1;
      patterns[103] = 12'b0_1_1_0_0_1_1_1_0_1_0_0;
      patterns[104] = 12'b0_1_1_0_1_0_0_0_1_0_1_1;
      patterns[105] = 12'b0_1_1_0_1_0_0_1_1_0_1_0;
      patterns[106] = 12'b0_1_1_0_1_0_1_0_1_0_0_1;
      patterns[107] = 12'b0_1_1_0_1_0_1_1_1_0_0_0;
      patterns[108] = 12'b0_1_1_0_1_1_0_0_0_1_1_1;
      patterns[109] = 12'b0_1_1_0_1_1_0_1_0_1_1_0;
      patterns[110] = 12'b0_1_1_0_1_1_1_0_0_1_0_1;
      patterns[111] = 12'b0_1_1_0_1_1_1_1_0_1_0_0;
      patterns[112] = 12'b0_1_1_1_0_0_0_0_0_1_1_1;
      patterns[113] = 12'b0_1_1_1_0_0_0_1_0_1_1_0;
      patterns[114] = 12'b0_1_1_1_0_0_1_0_0_1_0_1;
      patterns[115] = 12'b0_1_1_1_0_0_1_1_0_1_0_0;
      patterns[116] = 12'b0_1_1_1_0_1_0_0_0_0_1_1;
      patterns[117] = 12'b0_1_1_1_0_1_0_1_0_0_1_0;
      patterns[118] = 12'b0_1_1_1_0_1_1_0_0_0_0_1;
      patterns[119] = 12'b0_1_1_1_0_1_1_1_0_0_0_0;
      patterns[120] = 12'b0_1_1_1_1_0_0_0_1_1_1_1;
      patterns[121] = 12'b0_1_1_1_1_0_0_1_1_1_1_0;
      patterns[122] = 12'b0_1_1_1_1_0_1_0_1_1_0_1;
      patterns[123] = 12'b0_1_1_1_1_0_1_1_1_1_0_0;
      patterns[124] = 12'b0_1_1_1_1_1_0_0_1_0_1_1;
      patterns[125] = 12'b0_1_1_1_1_1_0_1_1_0_1_0;
      patterns[126] = 12'b0_1_1_1_1_1_1_0_1_0_0_1;
      patterns[127] = 12'b0_1_1_1_1_1_1_1_1_0_0_0;
      patterns[128] = 12'b1_0_0_0_0_0_0_0_1_0_0_0;
      patterns[129] = 12'b1_0_0_0_0_0_0_1_1_0_0_1;
      patterns[130] = 12'b1_0_0_0_0_0_1_0_1_0_1_0;
      patterns[131] = 12'b1_0_0_0_0_0_1_1_1_0_1_1;
      patterns[132] = 12'b1_0_0_0_0_1_0_0_1_1_0_0;
      patterns[133] = 12'b1_0_0_0_0_1_0_1_1_1_0_1;
      patterns[134] = 12'b1_0_0_0_0_1_1_0_1_1_1_0;
      patterns[135] = 12'b1_0_0_0_0_1_1_1_1_1_1_1;
      patterns[136] = 12'b1_0_0_0_1_0_0_0_0_0_0_0;
      patterns[137] = 12'b1_0_0_0_1_0_0_1_0_0_0_1;
      patterns[138] = 12'b1_0_0_0_1_0_1_0_0_0_1_0;
      patterns[139] = 12'b1_0_0_0_1_0_1_1_0_0_1_1;
      patterns[140] = 12'b1_0_0_0_1_1_0_0_0_1_0_0;
      patterns[141] = 12'b1_0_0_0_1_1_0_1_0_1_0_1;
      patterns[142] = 12'b1_0_0_0_1_1_1_0_0_1_1_0;
      patterns[143] = 12'b1_0_0_0_1_1_1_1_0_1_1_1;
      patterns[144] = 12'b1_0_0_1_0_0_0_0_0_1_0_0;
      patterns[145] = 12'b1_0_0_1_0_0_0_1_0_1_0_1;
      patterns[146] = 12'b1_0_0_1_0_0_1_0_0_1_1_0;
      patterns[147] = 12'b1_0_0_1_0_0_1_1_0_1_1_1;
      patterns[148] = 12'b1_0_0_1_0_1_0_0_1_0_0_0;
      patterns[149] = 12'b1_0_0_1_0_1_0_1_1_0_0_1;
      patterns[150] = 12'b1_0_0_1_0_1_1_0_1_0_1_0;
      patterns[151] = 12'b1_0_0_1_0_1_1_1_1_0_1_1;
      patterns[152] = 12'b1_0_0_1_1_0_0_0_0_1_0_0;
      patterns[153] = 12'b1_0_0_1_1_0_0_1_0_0_1_1;
      patterns[154] = 12'b1_0_0_1_1_0_1_0_0_0_1_0;
      patterns[155] = 12'b1_0_0_1_1_0_1_1_0_0_0_1;
      patterns[156] = 12'b1_0_0_1_1_1_0_0_0_0_0_0;
      patterns[157] = 12'b1_0_0_1_1_1_0_1_0_0_0_1;
      patterns[158] = 12'b1_0_0_1_1_1_1_0_0_0_1_0;
      patterns[159] = 12'b1_0_0_1_1_1_1_1_0_0_1_1;
      patterns[160] = 12'b1_0_1_0_0_0_0_0_0_1_1_0;
      patterns[161] = 12'b1_0_1_0_0_0_0_1_0_1_1_1;
      patterns[162] = 12'b1_0_1_0_0_0_1_0_1_0_0_0;
      patterns[163] = 12'b1_0_1_0_0_0_1_1_1_0_0_1;
      patterns[164] = 12'b1_0_1_0_0_1_0_0_1_0_1_0;
      patterns[165] = 12'b1_0_1_0_0_1_0_1_1_0_1_1;
      patterns[166] = 12'b1_0_1_0_0_1_1_0_1_1_0_0;
      patterns[167] = 12'b1_0_1_0_0_1_1_1_1_1_0_1;
      patterns[168] = 12'b1_0_1_0_1_0_0_0_0_0_1_0;
      patterns[169] = 12'b1_0_1_0_1_0_0_1_0_0_0_1;
      patterns[170] = 12'b1_0_1_0_1_0_1_0_0_0_0_0;
      patterns[171] = 12'b1_0_1_0_1_0_1_1_0_0_0_1;
      patterns[172] = 12'b1_0_1_0_1_1_0_0_0_0_1_0;
      patterns[173] = 12'b1_0_1_0_1_1_0_1_0_0_1_1;
      patterns[174] = 12'b1_0_1_0_1_1_1_0_0_1_0_0;
      patterns[175] = 12'b1_0_1_0_1_1_1_1_0_1_0_1;
      patterns[176] = 12'b1_0_1_1_0_0_0_0_0_0_1_0;
      patterns[177] = 12'b1_0_1_1_0_0_0_1_0_0_1_1;
      patterns[178] = 12'b1_0_1_1_0_0_1_0_0_1_0_0;
      patterns[179] = 12'b1_0_1_1_0_0_1_1_0_1_0_1;
      patterns[180] = 12'b1_0_1_1_0_1_0_0_0_1_1_0;
      patterns[181] = 12'b1_0_1_1_0_1_0_1_0_1_1_1;
      patterns[182] = 12'b1_0_1_1_0_1_1_0_1_0_0_0;
      patterns[183] = 12'b1_0_1_1_0_1_1_1_1_0_0_1;
      patterns[184] = 12'b1_0_1_1_1_0_0_0_0_1_1_0;
      patterns[185] = 12'b1_0_1_1_1_0_0_1_0_1_0_1;
      patterns[186] = 12'b1_0_1_1_1_0_1_0_0_1_0_0;
      patterns[187] = 12'b1_0_1_1_1_0_1_1_0_0_1_1;
      patterns[188] = 12'b1_0_1_1_1_1_0_0_0_0_1_0;
      patterns[189] = 12'b1_0_1_1_1_1_0_1_0_0_0_1;
      patterns[190] = 12'b1_0_1_1_1_1_1_0_0_0_0_0;
      patterns[191] = 12'b1_0_1_1_1_1_1_1_0_0_0_1;
      patterns[192] = 12'b1_1_0_0_0_0_0_0_0_1_1_1;
      patterns[193] = 12'b1_1_0_0_0_0_0_1_1_0_0_0;
      patterns[194] = 12'b1_1_0_0_0_0_1_0_1_0_0_1;
      patterns[195] = 12'b1_1_0_0_0_0_1_1_1_0_1_0;
      patterns[196] = 12'b1_1_0_0_0_1_0_0_1_0_1_1;
      patterns[197] = 12'b1_1_0_0_0_1_0_1_1_1_0_0;
      patterns[198] = 12'b1_1_0_0_0_1_1_0_1_1_0_1;
      patterns[199] = 12'b1_1_0_0_0_1_1_1_1_1_1_0;
      patterns[200] = 12'b1_1_0_0_1_0_0_0_0_0_0_1;
      patterns[201] = 12'b1_1_0_0_1_0_0_1_0_0_0_0;
      patterns[202] = 12'b1_1_0_0_1_0_1_0_0_0_0_1;
      patterns[203] = 12'b1_1_0_0_1_0_1_1_0_0_1_0;
      patterns[204] = 12'b1_1_0_0_1_1_0_0_0_0_1_1;
      patterns[205] = 12'b1_1_0_0_1_1_0_1_0_1_0_0;
      patterns[206] = 12'b1_1_0_0_1_1_1_0_0_1_0_1;
      patterns[207] = 12'b1_1_0_0_1_1_1_1_0_1_1_0;
      patterns[208] = 12'b1_1_0_1_0_0_0_0_0_0_1_1;
      patterns[209] = 12'b1_1_0_1_0_0_0_1_0_1_0_0;
      patterns[210] = 12'b1_1_0_1_0_0_1_0_0_1_0_1;
      patterns[211] = 12'b1_1_0_1_0_0_1_1_0_1_1_0;
      patterns[212] = 12'b1_1_0_1_0_1_0_0_0_1_1_1;
      patterns[213] = 12'b1_1_0_1_0_1_0_1_1_0_0_0;
      patterns[214] = 12'b1_1_0_1_0_1_1_0_1_0_0_1;
      patterns[215] = 12'b1_1_0_1_0_1_1_1_1_0_1_0;
      patterns[216] = 12'b1_1_0_1_1_0_0_0_0_1_0_1;
      patterns[217] = 12'b1_1_0_1_1_0_0_1_0_1_0_0;
      patterns[218] = 12'b1_1_0_1_1_0_1_0_0_0_1_1;
      patterns[219] = 12'b1_1_0_1_1_0_1_1_0_0_1_0;
      patterns[220] = 12'b1_1_0_1_1_1_0_0_0_0_0_1;
      patterns[221] = 12'b1_1_0_1_1_1_0_1_0_0_0_0;
      patterns[222] = 12'b1_1_0_1_1_1_1_0_0_0_0_1;
      patterns[223] = 12'b1_1_0_1_1_1_1_1_0_0_1_0;
      patterns[224] = 12'b1_1_1_0_0_0_0_0_0_1_0_1;
      patterns[225] = 12'b1_1_1_0_0_0_0_1_0_1_1_0;
      patterns[226] = 12'b1_1_1_0_0_0_1_0_0_1_1_1;
      patterns[227] = 12'b1_1_1_0_0_0_1_1_1_0_0_0;
      patterns[228] = 12'b1_1_1_0_0_1_0_0_1_0_0_1;
      patterns[229] = 12'b1_1_1_0_0_1_0_1_1_0_1_0;
      patterns[230] = 12'b1_1_1_0_0_1_1_0_1_0_1_1;
      patterns[231] = 12'b1_1_1_0_0_1_1_1_1_1_0_0;
      patterns[232] = 12'b1_1_1_0_1_0_0_0_0_0_1_1;
      patterns[233] = 12'b1_1_1_0_1_0_0_1_0_0_1_0;
      patterns[234] = 12'b1_1_1_0_1_0_1_0_0_0_0_1;
      patterns[235] = 12'b1_1_1_0_1_0_1_1_0_0_0_0;
      patterns[236] = 12'b1_1_1_0_1_1_0_0_0_0_0_1;
      patterns[237] = 12'b1_1_1_0_1_1_0_1_0_0_1_0;
      patterns[238] = 12'b1_1_1_0_1_1_1_0_0_0_1_1;
      patterns[239] = 12'b1_1_1_0_1_1_1_1_0_1_0_0;
      patterns[240] = 12'b1_1_1_1_0_0_0_0_0_0_0_1;
      patterns[241] = 12'b1_1_1_1_0_0_0_1_0_0_1_0;
      patterns[242] = 12'b1_1_1_1_0_0_1_0_0_0_1_1;
      patterns[243] = 12'b1_1_1_1_0_0_1_1_0_1_0_0;
      patterns[244] = 12'b1_1_1_1_0_1_0_0_0_1_0_1;
      patterns[245] = 12'b1_1_1_1_0_1_0_1_0_1_1_0;
      patterns[246] = 12'b1_1_1_1_0_1_1_0_0_1_1_1;
      patterns[247] = 12'b1_1_1_1_0_1_1_1_1_0_0_0;
      patterns[248] = 12'b1_1_1_1_1_0_0_0_0_1_1_1;
      patterns[249] = 12'b1_1_1_1_1_0_0_1_0_1_1_0;
      patterns[250] = 12'b1_1_1_1_1_0_1_0_0_1_0_1;
      patterns[251] = 12'b1_1_1_1_1_0_1_1_0_1_0_0;
      patterns[252] = 12'b1_1_1_1_1_1_0_0_0_0_1_1;
      patterns[253] = 12'b1_1_1_1_1_1_0_1_0_0_1_0;
      patterns[254] = 12'b1_1_1_1_1_1_1_0_0_0_0_1;
      patterns[255] = 12'b1_1_1_1_1_1_1_1_0_0_0_0;

      for (i = 0; i < 256; i = i + 1)
      begin
        B3 = patterns[i][11];
        A0 = patterns[i][10];
        A1 = patterns[i][9];
        A2 = patterns[i][8];
        A3 = patterns[i][7];
        B2 = patterns[i][6];
        B1 = patterns[i][5];
        B0 = patterns[i][4];
        #10;
        if (patterns[i][3] !== 1'hx)
        begin
          if (S3 !== patterns[i][3])
          begin
            $display("%d:S3: (assertion error). Expected %h, found %h", i, patterns[i][3], S3);
            $finish;
          end
        end
        if (patterns[i][2] !== 1'hx)
        begin
          if (S2 !== patterns[i][2])
          begin
            $display("%d:S2: (assertion error). Expected %h, found %h", i, patterns[i][2], S2);
            $finish;
          end
        end
        if (patterns[i][1] !== 1'hx)
        begin
          if (S1 !== patterns[i][1])
          begin
            $display("%d:S1: (assertion error). Expected %h, found %h", i, patterns[i][1], S1);
            $finish;
          end
        end
        if (patterns[i][0] !== 1'hx)
        begin
          if (S0 !== patterns[i][0])
          begin
            $display("%d:S0: (assertion error). Expected %h, found %h", i, patterns[i][0], S0);
            $finish;
          end
        end
      end

      $display("All tests passed.");
    end
  initial
  begin
    $dumpfile("SumadorRestador.vcd");
    $dumpvars(0, SumadorRestador_tb);
  end
    endmodule
